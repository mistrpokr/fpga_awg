module state_sel (
	state, out
);
	input state; 
	output out; 

	
endmodule