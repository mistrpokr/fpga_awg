module sin_table(input [9:0]address,
                 output reg[13:0]data);
    always @(*)
    begin
        case (address)
            10'd0: data    <= 14'd8192;
            10'd1: data    <= 14'd8242;
            10'd2: data    <= 14'd8292;
            10'd3: data    <= 14'd8342;
            10'd4: data    <= 14'd8393;
            10'd5: data    <= 14'd8443;
            10'd6: data    <= 14'd8493;
            10'd7: data    <= 14'd8543;
            10'd8: data    <= 14'd8593;
            10'd9: data    <= 14'd8644;
            10'd10: data   <= 14'd8694;
            10'd11: data   <= 14'd8744;
            10'd12: data   <= 14'd8794;
            10'd13: data   <= 14'd8844;
            10'd14: data   <= 14'd8894;
            10'd15: data   <= 14'd8944;
            10'd16: data   <= 14'd8994;
            10'd17: data   <= 14'd9044;
            10'd18: data   <= 14'd9094;
            10'd19: data   <= 14'd9144;
            10'd20: data   <= 14'd9194;
            10'd21: data   <= 14'd9244;
            10'd22: data   <= 14'd9294;
            10'd23: data   <= 14'd9344;
            10'd24: data   <= 14'd9394;
            10'd25: data   <= 14'd9443;
            10'd26: data   <= 14'd9493;
            10'd27: data   <= 14'd9542;
            10'd28: data   <= 14'd9592;
            10'd29: data   <= 14'd9642;
            10'd30: data   <= 14'd9691;
            10'd31: data   <= 14'd9740;
            10'd32: data   <= 14'd9790;
            10'd33: data   <= 14'd9839;
            10'd34: data   <= 14'd9888;
            10'd35: data   <= 14'd9937;
            10'd36: data   <= 14'd9986;
            10'd37: data   <= 14'd10035;
            10'd38: data   <= 14'd10084;
            10'd39: data   <= 14'd10133;
            10'd40: data   <= 14'd10182;
            10'd41: data   <= 14'd10231;
            10'd42: data   <= 14'd10279;
            10'd43: data   <= 14'd10328;
            10'd44: data   <= 14'd10376;
            10'd45: data   <= 14'd10425;
            10'd46: data   <= 14'd10473;
            10'd47: data   <= 14'd10521;
            10'd48: data   <= 14'd10570;
            10'd49: data   <= 14'd10618;
            10'd50: data   <= 14'd10666;
            10'd51: data   <= 14'd10713;
            10'd52: data   <= 14'd10761;
            10'd53: data   <= 14'd10809;
            10'd54: data   <= 14'd10856;
            10'd55: data   <= 14'd10904;
            10'd56: data   <= 14'd10951;
            10'd57: data   <= 14'd10999;
            10'd58: data   <= 14'd11046;
            10'd59: data   <= 14'd11093;
            10'd60: data   <= 14'd11140;
            10'd61: data   <= 14'd11187;
            10'd62: data   <= 14'd11233;
            10'd63: data   <= 14'd11280;
            10'd64: data   <= 14'd11326;
            10'd65: data   <= 14'd11373;
            10'd66: data   <= 14'd11419;
            10'd67: data   <= 14'd11465;
            10'd68: data   <= 14'd11511;
            10'd69: data   <= 14'd11557;
            10'd70: data   <= 14'd11603;
            10'd71: data   <= 14'd11649;
            10'd72: data   <= 14'd11694;
            10'd73: data   <= 14'd11739;
            10'd74: data   <= 14'd11785;
            10'd75: data   <= 14'd11830;
            10'd76: data   <= 14'd11875;
            10'd77: data   <= 14'd11920;
            10'd78: data   <= 14'd11964;
            10'd79: data   <= 14'd12009;
            10'd80: data   <= 14'd12053;
            10'd81: data   <= 14'd12097;
            10'd82: data   <= 14'd12142;
            10'd83: data   <= 14'd12186;
            10'd84: data   <= 14'd12229;
            10'd85: data   <= 14'd12273;
            10'd86: data   <= 14'd12316;
            10'd87: data   <= 14'd12360;
            10'd88: data   <= 14'd12403;
            10'd89: data   <= 14'd12446;
            10'd90: data   <= 14'd12489;
            10'd91: data   <= 14'd12532;
            10'd92: data   <= 14'd12574;
            10'd93: data   <= 14'd12617;
            10'd94: data   <= 14'd12659;
            10'd95: data   <= 14'd12701;
            10'd96: data   <= 14'd12743;
            10'd97: data   <= 14'd12784;
            10'd98: data   <= 14'd12826;
            10'd99: data   <= 14'd12867;
            10'd100: data  <= 14'd12909;
            10'd101: data  <= 14'd12950;
            10'd102: data  <= 14'd12990;
            10'd103: data  <= 14'd13031;
            10'd104: data  <= 14'd13071;
            10'd105: data  <= 14'd13112;
            10'd106: data  <= 14'd13152;
            10'd107: data  <= 14'd13192;
            10'd108: data  <= 14'd13231;
            10'd109: data  <= 14'd13271;
            10'd110: data  <= 14'd13310;
            10'd111: data  <= 14'd13349;
            10'd112: data  <= 14'd13388;
            10'd113: data  <= 14'd13427;
            10'd114: data  <= 14'd13466;
            10'd115: data  <= 14'd13504;
            10'd116: data  <= 14'd13542;
            10'd117: data  <= 14'd13580;
            10'd118: data  <= 14'd13618;
            10'd119: data  <= 14'd13656;
            10'd120: data  <= 14'd13693;
            10'd121: data  <= 14'd13730;
            10'd122: data  <= 14'd13767;
            10'd123: data  <= 14'd13804;
            10'd124: data  <= 14'd13840;
            10'd125: data  <= 14'd13877;
            10'd126: data  <= 14'd13913;
            10'd127: data  <= 14'd13948;
            10'd128: data  <= 14'd13984;
            10'd129: data  <= 14'd14020;
            10'd130: data  <= 14'd14055;
            10'd131: data  <= 14'd14090;
            10'd132: data  <= 14'd14125;
            10'd133: data  <= 14'd14159;
            10'd134: data  <= 14'd14193;
            10'd135: data  <= 14'd14228;
            10'd136: data  <= 14'd14261;
            10'd137: data  <= 14'd14295;
            10'd138: data  <= 14'd14328;
            10'd139: data  <= 14'd14362;
            10'd140: data  <= 14'd14395;
            10'd141: data  <= 14'd14427;
            10'd142: data  <= 14'd14460;
            10'd143: data  <= 14'd14492;
            10'd144: data  <= 14'd14524;
            10'd145: data  <= 14'd14556;
            10'd146: data  <= 14'd14587;
            10'd147: data  <= 14'd14619;
            10'd148: data  <= 14'd14650;
            10'd149: data  <= 14'd14680;
            10'd150: data  <= 14'd14711;
            10'd151: data  <= 14'd14741;
            10'd152: data  <= 14'd14771;
            10'd153: data  <= 14'd14801;
            10'd154: data  <= 14'd14831;
            10'd155: data  <= 14'd14860;
            10'd156: data  <= 14'd14889;
            10'd157: data  <= 14'd14918;
            10'd158: data  <= 14'd14947;
            10'd159: data  <= 14'd14975;
            10'd160: data  <= 14'd15003;
            10'd161: data  <= 14'd15031;
            10'd162: data  <= 14'd15058;
            10'd163: data  <= 14'd15086;
            10'd164: data  <= 14'd15113;
            10'd165: data  <= 14'd15139;
            10'd166: data  <= 14'd15166;
            10'd167: data  <= 14'd15192;
            10'd168: data  <= 14'd15218;
            10'd169: data  <= 14'd15244;
            10'd170: data  <= 14'd15269;
            10'd171: data  <= 14'd15294;
            10'd172: data  <= 14'd15319;
            10'd173: data  <= 14'd15344;
            10'd174: data  <= 14'd15368;
            10'd175: data  <= 14'd15392;
            10'd176: data  <= 14'd15416;
            10'd177: data  <= 14'd15440;
            10'd178: data  <= 14'd15463;
            10'd179: data  <= 14'd15486;
            10'd180: data  <= 14'd15509;
            10'd181: data  <= 14'd15531;
            10'd182: data  <= 14'd15553;
            10'd183: data  <= 14'd15575;
            10'd184: data  <= 14'd15597;
            10'd185: data  <= 14'd15618;
            10'd186: data  <= 14'd15639;
            10'd187: data  <= 14'd15660;
            10'd188: data  <= 14'd15681;
            10'd189: data  <= 14'd15701;
            10'd190: data  <= 14'd15721;
            10'd191: data  <= 14'd15741;
            10'd192: data  <= 14'd15760;
            10'd193: data  <= 14'd15779;
            10'd194: data  <= 14'd15798;
            10'd195: data  <= 14'd15816;
            10'd196: data  <= 14'd15835;
            10'd197: data  <= 14'd15853;
            10'd198: data  <= 14'd15870;
            10'd199: data  <= 14'd15888;
            10'd200: data  <= 14'd15905;
            10'd201: data  <= 14'd15921;
            10'd202: data  <= 14'd15938;
            10'd203: data  <= 14'd15954;
            10'd204: data  <= 14'd15970;
            10'd205: data  <= 14'd15986;
            10'd206: data  <= 14'd16001;
            10'd207: data  <= 14'd16016;
            10'd208: data  <= 14'd16031;
            10'd209: data  <= 14'd16045;
            10'd210: data  <= 14'd16059;
            10'd211: data  <= 14'd16073;
            10'd212: data  <= 14'd16087;
            10'd213: data  <= 14'd16100;
            10'd214: data  <= 14'd16113;
            10'd215: data  <= 14'd16126;
            10'd216: data  <= 14'd16138;
            10'd217: data  <= 14'd16150;
            10'd218: data  <= 14'd16162;
            10'd219: data  <= 14'd16173;
            10'd220: data  <= 14'd16184;
            10'd221: data  <= 14'd16195;
            10'd222: data  <= 14'd16206;
            10'd223: data  <= 14'd16216;
            10'd224: data  <= 14'd16226;
            10'd225: data  <= 14'd16236;
            10'd226: data  <= 14'd16245;
            10'd227: data  <= 14'd16254;
            10'd228: data  <= 14'd16263;
            10'd229: data  <= 14'd16271;
            10'd230: data  <= 14'd16279;
            10'd231: data  <= 14'd16287;
            10'd232: data  <= 14'd16295;
            10'd233: data  <= 14'd16302;
            10'd234: data  <= 14'd16309;
            10'd235: data  <= 14'd16316;
            10'd236: data  <= 14'd16322;
            10'd237: data  <= 14'd16328;
            10'd238: data  <= 14'd16334;
            10'd239: data  <= 14'd16339;
            10'd240: data  <= 14'd16344;
            10'd241: data  <= 14'd16349;
            10'd242: data  <= 14'd16353;
            10'd243: data  <= 14'd16357;
            10'd244: data  <= 14'd16361;
            10'd245: data  <= 14'd16365;
            10'd246: data  <= 14'd16368;
            10'd247: data  <= 14'd16371;
            10'd248: data  <= 14'd16374;
            10'd249: data  <= 14'd16376;
            10'd250: data  <= 14'd16378;
            10'd251: data  <= 14'd16380;
            10'd252: data  <= 14'd16381;
            10'd253: data  <= 14'd16382;
            10'd254: data  <= 14'd16383;
            10'd255: data  <= 14'd16383;
            10'd256: data  <= 14'd16384;
            10'd257: data  <= 14'd16383;
            10'd258: data  <= 14'd16383;
            10'd259: data  <= 14'd16382;
            10'd260: data  <= 14'd16381;
            10'd261: data  <= 14'd16380;
            10'd262: data  <= 14'd16378;
            10'd263: data  <= 14'd16376;
            10'd264: data  <= 14'd16374;
            10'd265: data  <= 14'd16371;
            10'd266: data  <= 14'd16368;
            10'd267: data  <= 14'd16365;
            10'd268: data  <= 14'd16361;
            10'd269: data  <= 14'd16357;
            10'd270: data  <= 14'd16353;
            10'd271: data  <= 14'd16349;
            10'd272: data  <= 14'd16344;
            10'd273: data  <= 14'd16339;
            10'd274: data  <= 14'd16334;
            10'd275: data  <= 14'd16328;
            10'd276: data  <= 14'd16322;
            10'd277: data  <= 14'd16316;
            10'd278: data  <= 14'd16309;
            10'd279: data  <= 14'd16302;
            10'd280: data  <= 14'd16295;
            10'd281: data  <= 14'd16287;
            10'd282: data  <= 14'd16279;
            10'd283: data  <= 14'd16271;
            10'd284: data  <= 14'd16263;
            10'd285: data  <= 14'd16254;
            10'd286: data  <= 14'd16245;
            10'd287: data  <= 14'd16236;
            10'd288: data  <= 14'd16226;
            10'd289: data  <= 14'd16216;
            10'd290: data  <= 14'd16206;
            10'd291: data  <= 14'd16195;
            10'd292: data  <= 14'd16184;
            10'd293: data  <= 14'd16173;
            10'd294: data  <= 14'd16162;
            10'd295: data  <= 14'd16150;
            10'd296: data  <= 14'd16138;
            10'd297: data  <= 14'd16126;
            10'd298: data  <= 14'd16113;
            10'd299: data  <= 14'd16100;
            10'd300: data  <= 14'd16087;
            10'd301: data  <= 14'd16073;
            10'd302: data  <= 14'd16059;
            10'd303: data  <= 14'd16045;
            10'd304: data  <= 14'd16031;
            10'd305: data  <= 14'd16016;
            10'd306: data  <= 14'd16001;
            10'd307: data  <= 14'd15986;
            10'd308: data  <= 14'd15970;
            10'd309: data  <= 14'd15954;
            10'd310: data  <= 14'd15938;
            10'd311: data  <= 14'd15921;
            10'd312: data  <= 14'd15905;
            10'd313: data  <= 14'd15888;
            10'd314: data  <= 14'd15870;
            10'd315: data  <= 14'd15853;
            10'd316: data  <= 14'd15835;
            10'd317: data  <= 14'd15816;
            10'd318: data  <= 14'd15798;
            10'd319: data  <= 14'd15779;
            10'd320: data  <= 14'd15760;
            10'd321: data  <= 14'd15741;
            10'd322: data  <= 14'd15721;
            10'd323: data  <= 14'd15701;
            10'd324: data  <= 14'd15681;
            10'd325: data  <= 14'd15660;
            10'd326: data  <= 14'd15639;
            10'd327: data  <= 14'd15618;
            10'd328: data  <= 14'd15597;
            10'd329: data  <= 14'd15575;
            10'd330: data  <= 14'd15553;
            10'd331: data  <= 14'd15531;
            10'd332: data  <= 14'd15509;
            10'd333: data  <= 14'd15486;
            10'd334: data  <= 14'd15463;
            10'd335: data  <= 14'd15440;
            10'd336: data  <= 14'd15416;
            10'd337: data  <= 14'd15392;
            10'd338: data  <= 14'd15368;
            10'd339: data  <= 14'd15344;
            10'd340: data  <= 14'd15319;
            10'd341: data  <= 14'd15294;
            10'd342: data  <= 14'd15269;
            10'd343: data  <= 14'd15244;
            10'd344: data  <= 14'd15218;
            10'd345: data  <= 14'd15192;
            10'd346: data  <= 14'd15166;
            10'd347: data  <= 14'd15139;
            10'd348: data  <= 14'd15113;
            10'd349: data  <= 14'd15086;
            10'd350: data  <= 14'd15058;
            10'd351: data  <= 14'd15031;
            10'd352: data  <= 14'd15003;
            10'd353: data  <= 14'd14975;
            10'd354: data  <= 14'd14947;
            10'd355: data  <= 14'd14918;
            10'd356: data  <= 14'd14889;
            10'd357: data  <= 14'd14860;
            10'd358: data  <= 14'd14831;
            10'd359: data  <= 14'd14801;
            10'd360: data  <= 14'd14771;
            10'd361: data  <= 14'd14741;
            10'd362: data  <= 14'd14711;
            10'd363: data  <= 14'd14680;
            10'd364: data  <= 14'd14650;
            10'd365: data  <= 14'd14619;
            10'd366: data  <= 14'd14587;
            10'd367: data  <= 14'd14556;
            10'd368: data  <= 14'd14524;
            10'd369: data  <= 14'd14492;
            10'd370: data  <= 14'd14460;
            10'd371: data  <= 14'd14427;
            10'd372: data  <= 14'd14395;
            10'd373: data  <= 14'd14362;
            10'd374: data  <= 14'd14328;
            10'd375: data  <= 14'd14295;
            10'd376: data  <= 14'd14261;
            10'd377: data  <= 14'd14228;
            10'd378: data  <= 14'd14193;
            10'd379: data  <= 14'd14159;
            10'd380: data  <= 14'd14125;
            10'd381: data  <= 14'd14090;
            10'd382: data  <= 14'd14055;
            10'd383: data  <= 14'd14020;
            10'd384: data  <= 14'd13984;
            10'd385: data  <= 14'd13948;
            10'd386: data  <= 14'd13913;
            10'd387: data  <= 14'd13877;
            10'd388: data  <= 14'd13840;
            10'd389: data  <= 14'd13804;
            10'd390: data  <= 14'd13767;
            10'd391: data  <= 14'd13730;
            10'd392: data  <= 14'd13693;
            10'd393: data  <= 14'd13656;
            10'd394: data  <= 14'd13618;
            10'd395: data  <= 14'd13580;
            10'd396: data  <= 14'd13542;
            10'd397: data  <= 14'd13504;
            10'd398: data  <= 14'd13466;
            10'd399: data  <= 14'd13427;
            10'd400: data  <= 14'd13388;
            10'd401: data  <= 14'd13349;
            10'd402: data  <= 14'd13310;
            10'd403: data  <= 14'd13271;
            10'd404: data  <= 14'd13231;
            10'd405: data  <= 14'd13192;
            10'd406: data  <= 14'd13152;
            10'd407: data  <= 14'd13112;
            10'd408: data  <= 14'd13071;
            10'd409: data  <= 14'd13031;
            10'd410: data  <= 14'd12990;
            10'd411: data  <= 14'd12950;
            10'd412: data  <= 14'd12909;
            10'd413: data  <= 14'd12867;
            10'd414: data  <= 14'd12826;
            10'd415: data  <= 14'd12784;
            10'd416: data  <= 14'd12743;
            10'd417: data  <= 14'd12701;
            10'd418: data  <= 14'd12659;
            10'd419: data  <= 14'd12617;
            10'd420: data  <= 14'd12574;
            10'd421: data  <= 14'd12532;
            10'd422: data  <= 14'd12489;
            10'd423: data  <= 14'd12446;
            10'd424: data  <= 14'd12403;
            10'd425: data  <= 14'd12360;
            10'd426: data  <= 14'd12316;
            10'd427: data  <= 14'd12273;
            10'd428: data  <= 14'd12229;
            10'd429: data  <= 14'd12186;
            10'd430: data  <= 14'd12142;
            10'd431: data  <= 14'd12097;
            10'd432: data  <= 14'd12053;
            10'd433: data  <= 14'd12009;
            10'd434: data  <= 14'd11964;
            10'd435: data  <= 14'd11920;
            10'd436: data  <= 14'd11875;
            10'd437: data  <= 14'd11830;
            10'd438: data  <= 14'd11785;
            10'd439: data  <= 14'd11739;
            10'd440: data  <= 14'd11694;
            10'd441: data  <= 14'd11649;
            10'd442: data  <= 14'd11603;
            10'd443: data  <= 14'd11557;
            10'd444: data  <= 14'd11511;
            10'd445: data  <= 14'd11465;
            10'd446: data  <= 14'd11419;
            10'd447: data  <= 14'd11373;
            10'd448: data  <= 14'd11326;
            10'd449: data  <= 14'd11280;
            10'd450: data  <= 14'd11233;
            10'd451: data  <= 14'd11187;
            10'd452: data  <= 14'd11140;
            10'd453: data  <= 14'd11093;
            10'd454: data  <= 14'd11046;
            10'd455: data  <= 14'd10999;
            10'd456: data  <= 14'd10951;
            10'd457: data  <= 14'd10904;
            10'd458: data  <= 14'd10856;
            10'd459: data  <= 14'd10809;
            10'd460: data  <= 14'd10761;
            10'd461: data  <= 14'd10713;
            10'd462: data  <= 14'd10666;
            10'd463: data  <= 14'd10618;
            10'd464: data  <= 14'd10570;
            10'd465: data  <= 14'd10521;
            10'd466: data  <= 14'd10473;
            10'd467: data  <= 14'd10425;
            10'd468: data  <= 14'd10376;
            10'd469: data  <= 14'd10328;
            10'd470: data  <= 14'd10279;
            10'd471: data  <= 14'd10231;
            10'd472: data  <= 14'd10182;
            10'd473: data  <= 14'd10133;
            10'd474: data  <= 14'd10084;
            10'd475: data  <= 14'd10035;
            10'd476: data  <= 14'd9986;
            10'd477: data  <= 14'd9937;
            10'd478: data  <= 14'd9888;
            10'd479: data  <= 14'd9839;
            10'd480: data  <= 14'd9790;
            10'd481: data  <= 14'd9740;
            10'd482: data  <= 14'd9691;
            10'd483: data  <= 14'd9642;
            10'd484: data  <= 14'd9592;
            10'd485: data  <= 14'd9542;
            10'd486: data  <= 14'd9493;
            10'd487: data  <= 14'd9443;
            10'd488: data  <= 14'd9394;
            10'd489: data  <= 14'd9344;
            10'd490: data  <= 14'd9294;
            10'd491: data  <= 14'd9244;
            10'd492: data  <= 14'd9194;
            10'd493: data  <= 14'd9144;
            10'd494: data  <= 14'd9094;
            10'd495: data  <= 14'd9044;
            10'd496: data  <= 14'd8994;
            10'd497: data  <= 14'd8944;
            10'd498: data  <= 14'd8894;
            10'd499: data  <= 14'd8844;
            10'd500: data  <= 14'd8794;
            10'd501: data  <= 14'd8744;
            10'd502: data  <= 14'd8694;
            10'd503: data  <= 14'd8644;
            10'd504: data  <= 14'd8593;
            10'd505: data  <= 14'd8543;
            10'd506: data  <= 14'd8493;
            10'd507: data  <= 14'd8443;
            10'd508: data  <= 14'd8393;
            10'd509: data  <= 14'd8342;
            10'd510: data  <= 14'd8292;
            10'd511: data  <= 14'd8242;
            10'd512: data  <= 14'd8192;
            10'd513: data  <= 14'd8141;
            10'd514: data  <= 14'd8091;
            10'd515: data  <= 14'd8041;
            10'd516: data  <= 14'd7990;
            10'd517: data  <= 14'd7940;
            10'd518: data  <= 14'd7890;
            10'd519: data  <= 14'd7840;
            10'd520: data  <= 14'd7790;
            10'd521: data  <= 14'd7739;
            10'd522: data  <= 14'd7689;
            10'd523: data  <= 14'd7639;
            10'd524: data  <= 14'd7589;
            10'd525: data  <= 14'd7539;
            10'd526: data  <= 14'd7489;
            10'd527: data  <= 14'd7439;
            10'd528: data  <= 14'd7389;
            10'd529: data  <= 14'd7339;
            10'd530: data  <= 14'd7289;
            10'd531: data  <= 14'd7239;
            10'd532: data  <= 14'd7189;
            10'd533: data  <= 14'd7139;
            10'd534: data  <= 14'd7089;
            10'd535: data  <= 14'd7039;
            10'd536: data  <= 14'd6989;
            10'd537: data  <= 14'd6940;
            10'd538: data  <= 14'd6890;
            10'd539: data  <= 14'd6841;
            10'd540: data  <= 14'd6791;
            10'd541: data  <= 14'd6741;
            10'd542: data  <= 14'd6692;
            10'd543: data  <= 14'd6643;
            10'd544: data  <= 14'd6593;
            10'd545: data  <= 14'd6544;
            10'd546: data  <= 14'd6495;
            10'd547: data  <= 14'd6446;
            10'd548: data  <= 14'd6397;
            10'd549: data  <= 14'd6348;
            10'd550: data  <= 14'd6299;
            10'd551: data  <= 14'd6250;
            10'd552: data  <= 14'd6201;
            10'd553: data  <= 14'd6152;
            10'd554: data  <= 14'd6104;
            10'd555: data  <= 14'd6055;
            10'd556: data  <= 14'd6007;
            10'd557: data  <= 14'd5958;
            10'd558: data  <= 14'd5910;
            10'd559: data  <= 14'd5862;
            10'd560: data  <= 14'd5813;
            10'd561: data  <= 14'd5765;
            10'd562: data  <= 14'd5717;
            10'd563: data  <= 14'd5670;
            10'd564: data  <= 14'd5622;
            10'd565: data  <= 14'd5574;
            10'd566: data  <= 14'd5527;
            10'd567: data  <= 14'd5479;
            10'd568: data  <= 14'd5432;
            10'd569: data  <= 14'd5384;
            10'd570: data  <= 14'd5337;
            10'd571: data  <= 14'd5290;
            10'd572: data  <= 14'd5243;
            10'd573: data  <= 14'd5196;
            10'd574: data  <= 14'd5150;
            10'd575: data  <= 14'd5103;
            10'd576: data  <= 14'd5057;
            10'd577: data  <= 14'd5010;
            10'd578: data  <= 14'd4964;
            10'd579: data  <= 14'd4918;
            10'd580: data  <= 14'd4872;
            10'd581: data  <= 14'd4826;
            10'd582: data  <= 14'd4780;
            10'd583: data  <= 14'd4734;
            10'd584: data  <= 14'd4689;
            10'd585: data  <= 14'd4644;
            10'd586: data  <= 14'd4598;
            10'd587: data  <= 14'd4553;
            10'd588: data  <= 14'd4508;
            10'd589: data  <= 14'd4463;
            10'd590: data  <= 14'd4419;
            10'd591: data  <= 14'd4374;
            10'd592: data  <= 14'd4330;
            10'd593: data  <= 14'd4286;
            10'd594: data  <= 14'd4241;
            10'd595: data  <= 14'd4197;
            10'd596: data  <= 14'd4154;
            10'd597: data  <= 14'd4110;
            10'd598: data  <= 14'd4067;
            10'd599: data  <= 14'd4023;
            10'd600: data  <= 14'd3980;
            10'd601: data  <= 14'd3937;
            10'd602: data  <= 14'd3894;
            10'd603: data  <= 14'd3851;
            10'd604: data  <= 14'd3809;
            10'd605: data  <= 14'd3766;
            10'd606: data  <= 14'd3724;
            10'd607: data  <= 14'd3682;
            10'd608: data  <= 14'd3640;
            10'd609: data  <= 14'd3599;
            10'd610: data  <= 14'd3557;
            10'd611: data  <= 14'd3516;
            10'd612: data  <= 14'd3474;
            10'd613: data  <= 14'd3433;
            10'd614: data  <= 14'd3393;
            10'd615: data  <= 14'd3352;
            10'd616: data  <= 14'd3312;
            10'd617: data  <= 14'd3271;
            10'd618: data  <= 14'd3231;
            10'd619: data  <= 14'd3191;
            10'd620: data  <= 14'd3152;
            10'd621: data  <= 14'd3112;
            10'd622: data  <= 14'd3073;
            10'd623: data  <= 14'd3034;
            10'd624: data  <= 14'd2995;
            10'd625: data  <= 14'd2956;
            10'd626: data  <= 14'd2917;
            10'd627: data  <= 14'd2879;
            10'd628: data  <= 14'd2841;
            10'd629: data  <= 14'd2803;
            10'd630: data  <= 14'd2765;
            10'd631: data  <= 14'd2727;
            10'd632: data  <= 14'd2690;
            10'd633: data  <= 14'd2653;
            10'd634: data  <= 14'd2616;
            10'd635: data  <= 14'd2579;
            10'd636: data  <= 14'd2543;
            10'd637: data  <= 14'd2506;
            10'd638: data  <= 14'd2470;
            10'd639: data  <= 14'd2435;
            10'd640: data  <= 14'd2399;
            10'd641: data  <= 14'd2363;
            10'd642: data  <= 14'd2328;
            10'd643: data  <= 14'd2293;
            10'd644: data  <= 14'd2258;
            10'd645: data  <= 14'd2224;
            10'd646: data  <= 14'd2190;
            10'd647: data  <= 14'd2155;
            10'd648: data  <= 14'd2122;
            10'd649: data  <= 14'd2088;
            10'd650: data  <= 14'd2055;
            10'd651: data  <= 14'd2021;
            10'd652: data  <= 14'd1988;
            10'd653: data  <= 14'd1956;
            10'd654: data  <= 14'd1923;
            10'd655: data  <= 14'd1891;
            10'd656: data  <= 14'd1859;
            10'd657: data  <= 14'd1827;
            10'd658: data  <= 14'd1796;
            10'd659: data  <= 14'd1764;
            10'd660: data  <= 14'd1733;
            10'd661: data  <= 14'd1703;
            10'd662: data  <= 14'd1672;
            10'd663: data  <= 14'd1642;
            10'd664: data  <= 14'd1612;
            10'd665: data  <= 14'd1582;
            10'd666: data  <= 14'd1552;
            10'd667: data  <= 14'd1523;
            10'd668: data  <= 14'd1494;
            10'd669: data  <= 14'd1465;
            10'd670: data  <= 14'd1436;
            10'd671: data  <= 14'd1408;
            10'd672: data  <= 14'd1380;
            10'd673: data  <= 14'd1352;
            10'd674: data  <= 14'd1325;
            10'd675: data  <= 14'd1297;
            10'd676: data  <= 14'd1270;
            10'd677: data  <= 14'd1244;
            10'd678: data  <= 14'd1217;
            10'd679: data  <= 14'd1191;
            10'd680: data  <= 14'd1165;
            10'd681: data  <= 14'd1139;
            10'd682: data  <= 14'd1114;
            10'd683: data  <= 14'd1089;
            10'd684: data  <= 14'd1064;
            10'd685: data  <= 14'd1039;
            10'd686: data  <= 14'd1015;
            10'd687: data  <= 14'd991;
            10'd688: data  <= 14'd967;
            10'd689: data  <= 14'd943;
            10'd690: data  <= 14'd920;
            10'd691: data  <= 14'd897;
            10'd692: data  <= 14'd874;
            10'd693: data  <= 14'd852;
            10'd694: data  <= 14'd830;
            10'd695: data  <= 14'd808;
            10'd696: data  <= 14'd786;
            10'd697: data  <= 14'd765;
            10'd698: data  <= 14'd744;
            10'd699: data  <= 14'd723;
            10'd700: data  <= 14'd702;
            10'd701: data  <= 14'd682;
            10'd702: data  <= 14'd662;
            10'd703: data  <= 14'd642;
            10'd704: data  <= 14'd623;
            10'd705: data  <= 14'd604;
            10'd706: data  <= 14'd585;
            10'd707: data  <= 14'd567;
            10'd708: data  <= 14'd548;
            10'd709: data  <= 14'd530;
            10'd710: data  <= 14'd513;
            10'd711: data  <= 14'd495;
            10'd712: data  <= 14'd478;
            10'd713: data  <= 14'd462;
            10'd714: data  <= 14'd445;
            10'd715: data  <= 14'd429;
            10'd716: data  <= 14'd413;
            10'd717: data  <= 14'd397;
            10'd718: data  <= 14'd382;
            10'd719: data  <= 14'd367;
            10'd720: data  <= 14'd352;
            10'd721: data  <= 14'd338;
            10'd722: data  <= 14'd324;
            10'd723: data  <= 14'd310;
            10'd724: data  <= 14'd296;
            10'd725: data  <= 14'd283;
            10'd726: data  <= 14'd270;
            10'd727: data  <= 14'd257;
            10'd728: data  <= 14'd245;
            10'd729: data  <= 14'd233;
            10'd730: data  <= 14'd221;
            10'd731: data  <= 14'd210;
            10'd732: data  <= 14'd199;
            10'd733: data  <= 14'd188;
            10'd734: data  <= 14'd177;
            10'd735: data  <= 14'd167;
            10'd736: data  <= 14'd157;
            10'd737: data  <= 14'd147;
            10'd738: data  <= 14'd138;
            10'd739: data  <= 14'd129;
            10'd740: data  <= 14'd120;
            10'd741: data  <= 14'd112;
            10'd742: data  <= 14'd104;
            10'd743: data  <= 14'd96;
            10'd744: data  <= 14'd88;
            10'd745: data  <= 14'd81;
            10'd746: data  <= 14'd74;
            10'd747: data  <= 14'd67;
            10'd748: data  <= 14'd61;
            10'd749: data  <= 14'd55;
            10'd750: data  <= 14'd49;
            10'd751: data  <= 14'd44;
            10'd752: data  <= 14'd39;
            10'd753: data  <= 14'd34;
            10'd754: data  <= 14'd30;
            10'd755: data  <= 14'd26;
            10'd756: data  <= 14'd22;
            10'd757: data  <= 14'd18;
            10'd758: data  <= 14'd15;
            10'd759: data  <= 14'd12;
            10'd760: data  <= 14'd9;
            10'd761: data  <= 14'd7;
            10'd762: data  <= 14'd5;
            10'd763: data  <= 14'd3;
            10'd764: data  <= 14'd2;
            10'd765: data  <= 14'd1;
            10'd766: data  <= 14'd0;
            10'd767: data  <= 14'd0;
            10'd768: data  <= 14'd0;
            10'd769: data  <= 14'd0;
            10'd770: data  <= 14'd0;
            10'd771: data  <= 14'd1;
            10'd772: data  <= 14'd2;
            10'd773: data  <= 14'd3;
            10'd774: data  <= 14'd5;
            10'd775: data  <= 14'd7;
            10'd776: data  <= 14'd9;
            10'd777: data  <= 14'd12;
            10'd778: data  <= 14'd15;
            10'd779: data  <= 14'd18;
            10'd780: data  <= 14'd22;
            10'd781: data  <= 14'd26;
            10'd782: data  <= 14'd30;
            10'd783: data  <= 14'd34;
            10'd784: data  <= 14'd39;
            10'd785: data  <= 14'd44;
            10'd786: data  <= 14'd49;
            10'd787: data  <= 14'd55;
            10'd788: data  <= 14'd61;
            10'd789: data  <= 14'd67;
            10'd790: data  <= 14'd74;
            10'd791: data  <= 14'd81;
            10'd792: data  <= 14'd88;
            10'd793: data  <= 14'd96;
            10'd794: data  <= 14'd104;
            10'd795: data  <= 14'd112;
            10'd796: data  <= 14'd120;
            10'd797: data  <= 14'd129;
            10'd798: data  <= 14'd138;
            10'd799: data  <= 14'd147;
            10'd800: data  <= 14'd157;
            10'd801: data  <= 14'd167;
            10'd802: data  <= 14'd177;
            10'd803: data  <= 14'd188;
            10'd804: data  <= 14'd199;
            10'd805: data  <= 14'd210;
            10'd806: data  <= 14'd221;
            10'd807: data  <= 14'd233;
            10'd808: data  <= 14'd245;
            10'd809: data  <= 14'd257;
            10'd810: data  <= 14'd270;
            10'd811: data  <= 14'd283;
            10'd812: data  <= 14'd296;
            10'd813: data  <= 14'd310;
            10'd814: data  <= 14'd324;
            10'd815: data  <= 14'd338;
            10'd816: data  <= 14'd352;
            10'd817: data  <= 14'd367;
            10'd818: data  <= 14'd382;
            10'd819: data  <= 14'd397;
            10'd820: data  <= 14'd413;
            10'd821: data  <= 14'd429;
            10'd822: data  <= 14'd445;
            10'd823: data  <= 14'd462;
            10'd824: data  <= 14'd478;
            10'd825: data  <= 14'd495;
            10'd826: data  <= 14'd513;
            10'd827: data  <= 14'd530;
            10'd828: data  <= 14'd548;
            10'd829: data  <= 14'd567;
            10'd830: data  <= 14'd585;
            10'd831: data  <= 14'd604;
            10'd832: data  <= 14'd623;
            10'd833: data  <= 14'd642;
            10'd834: data  <= 14'd662;
            10'd835: data  <= 14'd682;
            10'd836: data  <= 14'd702;
            10'd837: data  <= 14'd723;
            10'd838: data  <= 14'd744;
            10'd839: data  <= 14'd765;
            10'd840: data  <= 14'd786;
            10'd841: data  <= 14'd808;
            10'd842: data  <= 14'd830;
            10'd843: data  <= 14'd852;
            10'd844: data  <= 14'd874;
            10'd845: data  <= 14'd897;
            10'd846: data  <= 14'd920;
            10'd847: data  <= 14'd943;
            10'd848: data  <= 14'd967;
            10'd849: data  <= 14'd991;
            10'd850: data  <= 14'd1015;
            10'd851: data  <= 14'd1039;
            10'd852: data  <= 14'd1064;
            10'd853: data  <= 14'd1089;
            10'd854: data  <= 14'd1114;
            10'd855: data  <= 14'd1139;
            10'd856: data  <= 14'd1165;
            10'd857: data  <= 14'd1191;
            10'd858: data  <= 14'd1217;
            10'd859: data  <= 14'd1244;
            10'd860: data  <= 14'd1270;
            10'd861: data  <= 14'd1297;
            10'd862: data  <= 14'd1325;
            10'd863: data  <= 14'd1352;
            10'd864: data  <= 14'd1380;
            10'd865: data  <= 14'd1408;
            10'd866: data  <= 14'd1436;
            10'd867: data  <= 14'd1465;
            10'd868: data  <= 14'd1494;
            10'd869: data  <= 14'd1523;
            10'd870: data  <= 14'd1552;
            10'd871: data  <= 14'd1582;
            10'd872: data  <= 14'd1612;
            10'd873: data  <= 14'd1642;
            10'd874: data  <= 14'd1672;
            10'd875: data  <= 14'd1703;
            10'd876: data  <= 14'd1733;
            10'd877: data  <= 14'd1764;
            10'd878: data  <= 14'd1796;
            10'd879: data  <= 14'd1827;
            10'd880: data  <= 14'd1859;
            10'd881: data  <= 14'd1891;
            10'd882: data  <= 14'd1923;
            10'd883: data  <= 14'd1956;
            10'd884: data  <= 14'd1988;
            10'd885: data  <= 14'd2021;
            10'd886: data  <= 14'd2055;
            10'd887: data  <= 14'd2088;
            10'd888: data  <= 14'd2122;
            10'd889: data  <= 14'd2155;
            10'd890: data  <= 14'd2190;
            10'd891: data  <= 14'd2224;
            10'd892: data  <= 14'd2258;
            10'd893: data  <= 14'd2293;
            10'd894: data  <= 14'd2328;
            10'd895: data  <= 14'd2363;
            10'd896: data  <= 14'd2399;
            10'd897: data  <= 14'd2435;
            10'd898: data  <= 14'd2470;
            10'd899: data  <= 14'd2506;
            10'd900: data  <= 14'd2543;
            10'd901: data  <= 14'd2579;
            10'd902: data  <= 14'd2616;
            10'd903: data  <= 14'd2653;
            10'd904: data  <= 14'd2690;
            10'd905: data  <= 14'd2727;
            10'd906: data  <= 14'd2765;
            10'd907: data  <= 14'd2803;
            10'd908: data  <= 14'd2841;
            10'd909: data  <= 14'd2879;
            10'd910: data  <= 14'd2917;
            10'd911: data  <= 14'd2956;
            10'd912: data  <= 14'd2995;
            10'd913: data  <= 14'd3034;
            10'd914: data  <= 14'd3073;
            10'd915: data  <= 14'd3112;
            10'd916: data  <= 14'd3152;
            10'd917: data  <= 14'd3191;
            10'd918: data  <= 14'd3231;
            10'd919: data  <= 14'd3271;
            10'd920: data  <= 14'd3312;
            10'd921: data  <= 14'd3352;
            10'd922: data  <= 14'd3393;
            10'd923: data  <= 14'd3433;
            10'd924: data  <= 14'd3474;
            10'd925: data  <= 14'd3516;
            10'd926: data  <= 14'd3557;
            10'd927: data  <= 14'd3599;
            10'd928: data  <= 14'd3640;
            10'd929: data  <= 14'd3682;
            10'd930: data  <= 14'd3724;
            10'd931: data  <= 14'd3766;
            10'd932: data  <= 14'd3809;
            10'd933: data  <= 14'd3851;
            10'd934: data  <= 14'd3894;
            10'd935: data  <= 14'd3937;
            10'd936: data  <= 14'd3980;
            10'd937: data  <= 14'd4023;
            10'd938: data  <= 14'd4067;
            10'd939: data  <= 14'd4110;
            10'd940: data  <= 14'd4154;
            10'd941: data  <= 14'd4197;
            10'd942: data  <= 14'd4241;
            10'd943: data  <= 14'd4286;
            10'd944: data  <= 14'd4330;
            10'd945: data  <= 14'd4374;
            10'd946: data  <= 14'd4419;
            10'd947: data  <= 14'd4463;
            10'd948: data  <= 14'd4508;
            10'd949: data  <= 14'd4553;
            10'd950: data  <= 14'd4598;
            10'd951: data  <= 14'd4644;
            10'd952: data  <= 14'd4689;
            10'd953: data  <= 14'd4734;
            10'd954: data  <= 14'd4780;
            10'd955: data  <= 14'd4826;
            10'd956: data  <= 14'd4872;
            10'd957: data  <= 14'd4918;
            10'd958: data  <= 14'd4964;
            10'd959: data  <= 14'd5010;
            10'd960: data  <= 14'd5057;
            10'd961: data  <= 14'd5103;
            10'd962: data  <= 14'd5150;
            10'd963: data  <= 14'd5196;
            10'd964: data  <= 14'd5243;
            10'd965: data  <= 14'd5290;
            10'd966: data  <= 14'd5337;
            10'd967: data  <= 14'd5384;
            10'd968: data  <= 14'd5432;
            10'd969: data  <= 14'd5479;
            10'd970: data  <= 14'd5527;
            10'd971: data  <= 14'd5574;
            10'd972: data  <= 14'd5622;
            10'd973: data  <= 14'd5670;
            10'd974: data  <= 14'd5717;
            10'd975: data  <= 14'd5765;
            10'd976: data  <= 14'd5813;
            10'd977: data  <= 14'd5862;
            10'd978: data  <= 14'd5910;
            10'd979: data  <= 14'd5958;
            10'd980: data  <= 14'd6007;
            10'd981: data  <= 14'd6055;
            10'd982: data  <= 14'd6104;
            10'd983: data  <= 14'd6152;
            10'd984: data  <= 14'd6201;
            10'd985: data  <= 14'd6250;
            10'd986: data  <= 14'd6299;
            10'd987: data  <= 14'd6348;
            10'd988: data  <= 14'd6397;
            10'd989: data  <= 14'd6446;
            10'd990: data  <= 14'd6495;
            10'd991: data  <= 14'd6544;
            10'd992: data  <= 14'd6593;
            10'd993: data  <= 14'd6643;
            10'd994: data  <= 14'd6692;
            10'd995: data  <= 14'd6741;
            10'd996: data  <= 14'd6791;
            10'd997: data  <= 14'd6841;
            10'd998: data  <= 14'd6890;
            10'd999: data  <= 14'd6940;
            10'd1000: data <= 14'd6989;
            10'd1001: data <= 14'd7039;
            10'd1002: data <= 14'd7089;
            10'd1003: data <= 14'd7139;
            10'd1004: data <= 14'd7189;
            10'd1005: data <= 14'd7239;
            10'd1006: data <= 14'd7289;
            10'd1007: data <= 14'd7339;
            10'd1008: data <= 14'd7389;
            10'd1009: data <= 14'd7439;
            10'd1010: data <= 14'd7489;
            10'd1011: data <= 14'd7539;
            10'd1012: data <= 14'd7589;
            10'd1013: data <= 14'd7639;
            10'd1014: data <= 14'd7689;
            10'd1015: data <= 14'd7739;
            10'd1016: data <= 14'd7790;
            10'd1017: data <= 14'd7840;
            10'd1018: data <= 14'd7890;
            10'd1019: data <= 14'd7940;
            10'd1020: data <= 14'd7990;
            10'd1021: data <= 14'd8041;
            10'd1022: data <= 14'd8091;
            10'd1023: data <= 14'd8141;
        endcase
    end
endmodule
