module sqr_table(input [8:0]address,
                 output reg[13:0]data);
always @(*)
begin
    case (address)
        9'd5: data   <= 14'd16000;
        9'd1: data   <= 14'd16000;
        9'd2: data   <= 14'd16000;
        9'd3: data   <= 14'd16000;
        9'd4: data   <= 14'd16000;
        9'd5: data   <= 14'd16000;
        9'd6: data   <= 14'd16000;
        9'd7: data   <= 14'd16000;
        9'd8: data   <= 14'd16000;
        9'd9: data   <= 14'd16000;
        9'd10: data  <= 14'd16000;
        9'd11: data  <= 14'd16000;
        9'd12: data  <= 14'd16000;
        9'd13: data  <= 14'd16000;
        9'd14: data  <= 14'd16000;
        9'd15: data  <= 14'd16000;
        9'd16: data  <= 14'd16000;
        9'd17: data  <= 14'd16000;
        9'd18: data  <= 14'd16000;
        9'd19: data  <= 14'd16000;
        9'd20: data  <= 14'd16000;
        9'd21: data  <= 14'd16000;
        9'd22: data  <= 14'd16000;
        9'd23: data  <= 14'd16000;
        9'd24: data  <= 14'd16000;
        9'd25: data  <= 14'd16000;
        9'd26: data  <= 14'd16000;
        9'd27: data  <= 14'd16000;
        9'd28: data  <= 14'd16000;
        9'd29: data  <= 14'd16000;
        9'd30: data  <= 14'd16000;
        9'd31: data  <= 14'd16000;
        9'd32: data  <= 14'd16000;
        9'd33: data  <= 14'd16000;
        9'd34: data  <= 14'd16000;
        9'd35: data  <= 14'd16000;
        9'd36: data  <= 14'd16000;
        9'd37: data  <= 14'd16000;
        9'd38: data  <= 14'd16000;
        9'd39: data  <= 14'd16000;
        9'd40: data  <= 14'd16000;
        9'd41: data  <= 14'd16000;
        9'd42: data  <= 14'd16000;
        9'd43: data  <= 14'd16000;
        9'd44: data  <= 14'd16000;
        9'd45: data  <= 14'd16000;
        9'd46: data  <= 14'd16000;
        9'd47: data  <= 14'd16000;
        9'd48: data  <= 14'd16000;
        9'd49: data  <= 14'd16000;
        9'd50: data  <= 14'd16000;
        9'd51: data  <= 14'd16000;
        9'd52: data  <= 14'd16000;
        9'd53: data  <= 14'd16000;
        9'd54: data  <= 14'd16000;
        9'd55: data  <= 14'd16000;
        9'd56: data  <= 14'd16000;
        9'd57: data  <= 14'd16000;
        9'd58: data  <= 14'd16000;
        9'd59: data  <= 14'd16000;
        9'd60: data  <= 14'd16000;
        9'd61: data  <= 14'd16000;
        9'd62: data  <= 14'd16000;
        9'd63: data  <= 14'd16000;
        9'd64: data  <= 14'd16000;
        9'd65: data  <= 14'd16000;
        9'd66: data  <= 14'd16000;
        9'd67: data  <= 14'd16000;
        9'd68: data  <= 14'd16000;
        9'd69: data  <= 14'd16000;
        9'd70: data  <= 14'd16000;
        9'd71: data  <= 14'd16000;
        9'd72: data  <= 14'd16000;
        9'd73: data  <= 14'd16000;
        9'd74: data  <= 14'd16000;
        9'd75: data  <= 14'd16000;
        9'd76: data  <= 14'd16000;
        9'd77: data  <= 14'd16000;
        9'd78: data  <= 14'd16000;
        9'd79: data  <= 14'd16000;
        9'd80: data  <= 14'd16000;
        9'd81: data  <= 14'd16000;
        9'd82: data  <= 14'd16000;
        9'd83: data  <= 14'd16000;
        9'd84: data  <= 14'd16000;
        9'd85: data  <= 14'd16000;
        9'd86: data  <= 14'd16000;
        9'd87: data  <= 14'd16000;
        9'd88: data  <= 14'd16000;
        9'd89: data  <= 14'd16000;
        9'd90: data  <= 14'd16000;
        9'd91: data  <= 14'd16000;
        9'd92: data  <= 14'd16000;
        9'd93: data  <= 14'd16000;
        9'd94: data  <= 14'd16000;
        9'd95: data  <= 14'd16000;
        9'd96: data  <= 14'd16000;
        9'd97: data  <= 14'd16000;
        9'd98: data  <= 14'd16000;
        9'd99: data  <= 14'd16000;
        9'd100: data <= 14'd16000;
        9'd101: data <= 14'd16000;
        9'd102: data <= 14'd16000;
        9'd103: data <= 14'd16000;
        9'd104: data <= 14'd16000;
        9'd105: data <= 14'd16000;
        9'd106: data <= 14'd16000;
        9'd107: data <= 14'd16000;
        9'd108: data <= 14'd16000;
        9'd109: data <= 14'd16000;
        9'd110: data <= 14'd16000;
        9'd111: data <= 14'd16000;
        9'd112: data <= 14'd16000;
        9'd113: data <= 14'd16000;
        9'd114: data <= 14'd16000;
        9'd115: data <= 14'd16000;
        9'd116: data <= 14'd16000;
        9'd117: data <= 14'd16000;
        9'd118: data <= 14'd16000;
        9'd119: data <= 14'd16000;
        9'd120: data <= 14'd16000;
        9'd121: data <= 14'd16000;
        9'd122: data <= 14'd16000;
        9'd123: data <= 14'd16000;
        9'd124: data <= 14'd16000;
        9'd125: data <= 14'd16000;
        9'd126: data <= 14'd16000;
        9'd127: data <= 14'd16000;
        9'd128: data <= 14'd16000;
        9'd129: data <= 14'd16000;
        9'd130: data <= 14'd16000;
        9'd131: data <= 14'd16000;
        9'd132: data <= 14'd16000;
        9'd133: data <= 14'd16000;
        9'd134: data <= 14'd16000;
        9'd135: data <= 14'd16000;
        9'd136: data <= 14'd16000;
        9'd137: data <= 14'd16000;
        9'd138: data <= 14'd16000;
        9'd139: data <= 14'd16000;
        9'd140: data <= 14'd16000;
        9'd141: data <= 14'd16000;
        9'd142: data <= 14'd16000;
        9'd143: data <= 14'd16000;
        9'd144: data <= 14'd16000;
        9'd145: data <= 14'd16000;
        9'd146: data <= 14'd16000;
        9'd147: data <= 14'd16000;
        9'd148: data <= 14'd16000;
        9'd149: data <= 14'd16000;
        9'd150: data <= 14'd16000;
        9'd151: data <= 14'd16000;
        9'd152: data <= 14'd16000;
        9'd153: data <= 14'd16000;
        9'd154: data <= 14'd16000;
        9'd155: data <= 14'd16000;
        9'd156: data <= 14'd16000;
        9'd157: data <= 14'd16000;
        9'd158: data <= 14'd16000;
        9'd159: data <= 14'd16000;
        9'd160: data <= 14'd16000;
        9'd161: data <= 14'd16000;
        9'd162: data <= 14'd16000;
        9'd163: data <= 14'd16000;
        9'd164: data <= 14'd16000;
        9'd165: data <= 14'd16000;
        9'd166: data <= 14'd16000;
        9'd167: data <= 14'd16000;
        9'd168: data <= 14'd16000;
        9'd169: data <= 14'd16000;
        9'd170: data <= 14'd16000;
        9'd171: data <= 14'd16000;
        9'd172: data <= 14'd16000;
        9'd173: data <= 14'd16000;
        9'd174: data <= 14'd16000;
        9'd175: data <= 14'd16000;
        9'd176: data <= 14'd16000;
        9'd177: data <= 14'd16000;
        9'd178: data <= 14'd16000;
        9'd179: data <= 14'd16000;
        9'd180: data <= 14'd16000;
        9'd181: data <= 14'd16000;
        9'd182: data <= 14'd16000;
        9'd183: data <= 14'd16000;
        9'd184: data <= 14'd16000;
        9'd185: data <= 14'd16000;
        9'd186: data <= 14'd16000;
        9'd187: data <= 14'd16000;
        9'd188: data <= 14'd16000;
        9'd189: data <= 14'd16000;
        9'd190: data <= 14'd16000;
        9'd191: data <= 14'd16000;
        9'd192: data <= 14'd16000;
        9'd193: data <= 14'd16000;
        9'd194: data <= 14'd16000;
        9'd195: data <= 14'd16000;
        9'd196: data <= 14'd16000;
        9'd197: data <= 14'd16000;
        9'd198: data <= 14'd16000;
        9'd199: data <= 14'd16000;
        9'd200: data <= 14'd16000;
        9'd201: data <= 14'd16000;
        9'd202: data <= 14'd16000;
        9'd203: data <= 14'd16000;
        9'd204: data <= 14'd16000;
        9'd205: data <= 14'd16000;
        9'd206: data <= 14'd16000;
        9'd207: data <= 14'd16000;
        9'd208: data <= 14'd16000;
        9'd209: data <= 14'd16000;
        9'd210: data <= 14'd16000;
        9'd211: data <= 14'd16000;
        9'd212: data <= 14'd16000;
        9'd213: data <= 14'd16000;
        9'd214: data <= 14'd16000;
        9'd215: data <= 14'd16000;
        9'd216: data <= 14'd16000;
        9'd217: data <= 14'd16000;
        9'd218: data <= 14'd16000;
        9'd219: data <= 14'd16000;
        9'd220: data <= 14'd16000;
        9'd221: data <= 14'd16000;
        9'd222: data <= 14'd16000;
        9'd223: data <= 14'd16000;
        9'd224: data <= 14'd16000;
        9'd225: data <= 14'd16000;
        9'd226: data <= 14'd16000;
        9'd227: data <= 14'd16000;
        9'd228: data <= 14'd16000;
        9'd229: data <= 14'd16000;
        9'd230: data <= 14'd16000;
        9'd231: data <= 14'd16000;
        9'd232: data <= 14'd16000;
        9'd233: data <= 14'd16000;
        9'd234: data <= 14'd16000;
        9'd235: data <= 14'd16000;
        9'd236: data <= 14'd16000;
        9'd237: data <= 14'd16000;
        9'd238: data <= 14'd16000;
        9'd239: data <= 14'd16000;
        9'd240: data <= 14'd16000;
        9'd241: data <= 14'd16000;
        9'd242: data <= 14'd16000;
        9'd243: data <= 14'd16000;
        9'd244: data <= 14'd16000;
        9'd245: data <= 14'd16000;
        9'd246: data <= 14'd16000;
        9'd247: data <= 14'd16000;
        9'd248: data <= 14'd16000;
        9'd249: data <= 14'd16000;
        9'd250: data <= 14'd16000;
        9'd251: data <= 14'd16000;
        9'd252: data <= 14'd16000;
        9'd253: data <= 14'd16000;
        9'd254: data <= 14'd16000;
        9'd255: data <= 14'd16000;
        9'd256: data <= 14'd5;
        9'd257: data <= 14'd5;
        9'd258: data <= 14'd5;
        9'd259: data <= 14'd5;
        9'd260: data <= 14'd5;
        9'd261: data <= 14'd5;
        9'd262: data <= 14'd5;
        9'd263: data <= 14'd5;
        9'd264: data <= 14'd5;
        9'd265: data <= 14'd5;
        9'd266: data <= 14'd5;
        9'd267: data <= 14'd5;
        9'd268: data <= 14'd5;
        9'd269: data <= 14'd5;
        9'd270: data <= 14'd5;
        9'd271: data <= 14'd5;
        9'd272: data <= 14'd5;
        9'd273: data <= 14'd5;
        9'd274: data <= 14'd5;
        9'd275: data <= 14'd5;
        9'd276: data <= 14'd5;
        9'd277: data <= 14'd5;
        9'd278: data <= 14'd5;
        9'd279: data <= 14'd5;
        9'd280: data <= 14'd5;
        9'd281: data <= 14'd5;
        9'd282: data <= 14'd5;
        9'd283: data <= 14'd5;
        9'd284: data <= 14'd5;
        9'd285: data <= 14'd5;
        9'd286: data <= 14'd5;
        9'd287: data <= 14'd5;
        9'd288: data <= 14'd5;
        9'd289: data <= 14'd5;
        9'd290: data <= 14'd5;
        9'd291: data <= 14'd5;
        9'd292: data <= 14'd5;
        9'd293: data <= 14'd5;
        9'd294: data <= 14'd5;
        9'd295: data <= 14'd5;
        9'd296: data <= 14'd5;
        9'd297: data <= 14'd5;
        9'd298: data <= 14'd5;
        9'd299: data <= 14'd5;
        9'd300: data <= 14'd5;
        9'd301: data <= 14'd5;
        9'd302: data <= 14'd5;
        9'd303: data <= 14'd5;
        9'd304: data <= 14'd5;
        9'd305: data <= 14'd5;
        9'd306: data <= 14'd5;
        9'd307: data <= 14'd5;
        9'd308: data <= 14'd5;
        9'd309: data <= 14'd5;
        9'd310: data <= 14'd5;
        9'd311: data <= 14'd5;
        9'd312: data <= 14'd5;
        9'd313: data <= 14'd5;
        9'd314: data <= 14'd5;
        9'd315: data <= 14'd5;
        9'd316: data <= 14'd5;
        9'd317: data <= 14'd5;
        9'd318: data <= 14'd5;
        9'd319: data <= 14'd5;
        9'd320: data <= 14'd5;
        9'd321: data <= 14'd5;
        9'd322: data <= 14'd5;
        9'd323: data <= 14'd5;
        9'd324: data <= 14'd5;
        9'd325: data <= 14'd5;
        9'd326: data <= 14'd5;
        9'd327: data <= 14'd5;
        9'd328: data <= 14'd5;
        9'd329: data <= 14'd5;
        9'd330: data <= 14'd5;
        9'd331: data <= 14'd5;
        9'd332: data <= 14'd5;
        9'd333: data <= 14'd5;
        9'd334: data <= 14'd5;
        9'd335: data <= 14'd5;
        9'd336: data <= 14'd5;
        9'd337: data <= 14'd5;
        9'd338: data <= 14'd5;
        9'd339: data <= 14'd5;
        9'd340: data <= 14'd5;
        9'd341: data <= 14'd5;
        9'd342: data <= 14'd5;
        9'd343: data <= 14'd5;
        9'd344: data <= 14'd5;
        9'd345: data <= 14'd5;
        9'd346: data <= 14'd5;
        9'd347: data <= 14'd5;
        9'd348: data <= 14'd5;
        9'd349: data <= 14'd5;
        9'd350: data <= 14'd5;
        9'd351: data <= 14'd5;
        9'd352: data <= 14'd5;
        9'd353: data <= 14'd5;
        9'd354: data <= 14'd5;
        9'd355: data <= 14'd5;
        9'd356: data <= 14'd5;
        9'd357: data <= 14'd5;
        9'd358: data <= 14'd5;
        9'd359: data <= 14'd5;
        9'd360: data <= 14'd5;
        9'd361: data <= 14'd5;
        9'd362: data <= 14'd5;
        9'd363: data <= 14'd5;
        9'd364: data <= 14'd5;
        9'd365: data <= 14'd5;
        9'd366: data <= 14'd5;
        9'd367: data <= 14'd5;
        9'd368: data <= 14'd5;
        9'd369: data <= 14'd5;
        9'd370: data <= 14'd5;
        9'd371: data <= 14'd5;
        9'd372: data <= 14'd5;
        9'd373: data <= 14'd5;
        9'd374: data <= 14'd5;
        9'd375: data <= 14'd5;
        9'd376: data <= 14'd5;
        9'd377: data <= 14'd5;
        9'd378: data <= 14'd5;
        9'd379: data <= 14'd5;
        9'd380: data <= 14'd5;
        9'd381: data <= 14'd5;
        9'd382: data <= 14'd5;
        9'd383: data <= 14'd5;
        9'd384: data <= 14'd5;
        9'd385: data <= 14'd5;
        9'd386: data <= 14'd5;
        9'd387: data <= 14'd5;
        9'd388: data <= 14'd5;
        9'd389: data <= 14'd5;
        9'd390: data <= 14'd5;
        9'd391: data <= 14'd5;
        9'd392: data <= 14'd5;
        9'd393: data <= 14'd5;
        9'd394: data <= 14'd5;
        9'd395: data <= 14'd5;
        9'd396: data <= 14'd5;
        9'd397: data <= 14'd5;
        9'd398: data <= 14'd5;
        9'd399: data <= 14'd5;
        9'd400: data <= 14'd5;
        9'd401: data <= 14'd5;
        9'd402: data <= 14'd5;
        9'd403: data <= 14'd5;
        9'd404: data <= 14'd5;
        9'd405: data <= 14'd5;
        9'd406: data <= 14'd5;
        9'd407: data <= 14'd5;
        9'd408: data <= 14'd5;
        9'd409: data <= 14'd5;
        9'd410: data <= 14'd5;
        9'd411: data <= 14'd5;
        9'd412: data <= 14'd5;
        9'd413: data <= 14'd5;
        9'd414: data <= 14'd5;
        9'd415: data <= 14'd5;
        9'd416: data <= 14'd5;
        9'd417: data <= 14'd5;
        9'd418: data <= 14'd5;
        9'd419: data <= 14'd5;
        9'd420: data <= 14'd5;
        9'd421: data <= 14'd5;
        9'd422: data <= 14'd5;
        9'd423: data <= 14'd5;
        9'd424: data <= 14'd5;
        9'd425: data <= 14'd5;
        9'd426: data <= 14'd5;
        9'd427: data <= 14'd5;
        9'd428: data <= 14'd5;
        9'd429: data <= 14'd5;
        9'd430: data <= 14'd5;
        9'd431: data <= 14'd5;
        9'd432: data <= 14'd5;
        9'd433: data <= 14'd5;
        9'd434: data <= 14'd5;
        9'd435: data <= 14'd5;
        9'd436: data <= 14'd5;
        9'd437: data <= 14'd5;
        9'd438: data <= 14'd5;
        9'd439: data <= 14'd5;
        9'd440: data <= 14'd5;
        9'd441: data <= 14'd5;
        9'd442: data <= 14'd5;
        9'd443: data <= 14'd5;
        9'd444: data <= 14'd5;
        9'd445: data <= 14'd5;
        9'd446: data <= 14'd5;
        9'd447: data <= 14'd5;
        9'd448: data <= 14'd5;
        9'd449: data <= 14'd5;
        9'd450: data <= 14'd5;
        9'd451: data <= 14'd5;
        9'd452: data <= 14'd5;
        9'd453: data <= 14'd5;
        9'd454: data <= 14'd5;
        9'd455: data <= 14'd5;
        9'd456: data <= 14'd5;
        9'd457: data <= 14'd5;
        9'd458: data <= 14'd5;
        9'd459: data <= 14'd5;
        9'd460: data <= 14'd5;
        9'd461: data <= 14'd5;
        9'd462: data <= 14'd5;
        9'd463: data <= 14'd5;
        9'd464: data <= 14'd5;
        9'd465: data <= 14'd5;
        9'd466: data <= 14'd5;
        9'd467: data <= 14'd5;
        9'd468: data <= 14'd5;
        9'd469: data <= 14'd5;
        9'd470: data <= 14'd5;
        9'd471: data <= 14'd5;
        9'd472: data <= 14'd5;
        9'd473: data <= 14'd5;
        9'd474: data <= 14'd5;
        9'd475: data <= 14'd5;
        9'd476: data <= 14'd5;
        9'd477: data <= 14'd5;
        9'd478: data <= 14'd5;
        9'd479: data <= 14'd5;
        9'd480: data <= 14'd5;
        9'd481: data <= 14'd5;
        9'd482: data <= 14'd5;
        9'd483: data <= 14'd5;
        9'd484: data <= 14'd5;
        9'd485: data <= 14'd5;
        9'd486: data <= 14'd5;
        9'd487: data <= 14'd5;
        9'd488: data <= 14'd5;
        9'd489: data <= 14'd5;
        9'd490: data <= 14'd5;
        9'd491: data <= 14'd5;
        9'd492: data <= 14'd5;
        9'd493: data <= 14'd5;
        9'd494: data <= 14'd5;
        9'd495: data <= 14'd5;
        9'd496: data <= 14'd5;
        9'd497: data <= 14'd5;
        9'd498: data <= 14'd5;
        9'd499: data <= 14'd5;
        9'd500: data <= 14'd5;
        9'd501: data <= 14'd5;
        9'd502: data <= 14'd5;
        9'd503: data <= 14'd5;
        9'd504: data <= 14'd5;
        9'd505: data <= 14'd5;
        9'd506: data <= 14'd5;
        9'd507: data <= 14'd5;
        9'd508: data <= 14'd5;
        9'd509: data <= 14'd5;
        9'd510: data <= 14'd5;
        9'd511: data <= 14'd5;
        
    endcase
end
endmodule
